1
7
2
3
example
_ _ _ _ _ _ _ 
EASY
